//------------------------------------------------------------------------
// MIPS-Subset Instructions
//------------------------------------------------------------------------

// load word
module LW
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// store word
module SW
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// jump
module J
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// jump register
module JR
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// jump and link
module JAL
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// branch on equal
module BEQ
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// branch on not equal
module BNE
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// bitwise exclusive OR immediate
module XORI
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// add immediate (with overflow)
module ADDI
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// add (with overflow)
module ADD
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// subtract
module SUB
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule


// set less than
module SLT
(
input 	    x,
output reg  y
);

    assign y = x;

endmodule
